/*Copyright 2020-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @23
module pa_fmau_lza_single(
  addend,
  lza_result,
  sub_vld,
  summand,
  upper_limit
);

// &Ports; @24
input   [52:0]  addend;      
input           sub_vld;     
input   [52:0]  summand;     
input   [52:0]  upper_limit; 
output  [6 :0]  lza_result;  

// &Regs; @25
reg     [6 :0]  lza_result;  

// &Wires; @26
wire    [52:0]  addend;      
wire    [52:0]  carry_d;     
wire    [52:0]  carry_g;     
wire    [52:0]  carry_p;     
wire    [52:0]  data_for_ff1; 
wire    [52:0]  lza_precod;  
wire            sub_vld;     
wire    [52:0]  summand;     
wire    [52:0]  upper_limit; 


parameter DATA_WIDTH = 53;
//==========================================================
//                   Signal Pre-encode
//==========================================================
//----------------------------------------------------------
//                   Signal preparation
//----------------------------------------------------------
// carry_p: carry propagete
// carry_g: carry generate
// carry_d: carry delete
assign carry_p[DATA_WIDTH-1:0] =   summand[DATA_WIDTH-1:0] ^ addend[DATA_WIDTH-1:0];
assign carry_g[DATA_WIDTH-1:0] =   summand[DATA_WIDTH-1:0] & addend[DATA_WIDTH-1:0];
assign carry_d[DATA_WIDTH-1:0] = ~(summand[DATA_WIDTH-1:0] | addend[DATA_WIDTH-1:0]);
//----------------------------------------------------------
//                   Signal decode
//----------------------------------------------------------
//pre-predecode for leading zero anticipation
assign lza_precod[0] = 
     carry_p[1] && (carry_g[0] && sub_vld || carry_d[0])
 || !carry_p[1] && (carry_d[0] && sub_vld || carry_g[0]);

assign lza_precod[DATA_WIDTH-1] = 
     sub_vld && (carry_g[DATA_WIDTH-1] && !carry_d[DATA_WIDTH-2] 
 ||  carry_d[DATA_WIDTH-1] && !carry_g[DATA_WIDTH-2])
 || !sub_vld && (carry_d[DATA_WIDTH-1] && !carry_d[DATA_WIDTH-2] 
 || !carry_d[DATA_WIDTH-1]);

assign lza_precod[DATA_WIDTH-2:1] = 
    carry_p[DATA_WIDTH-1:2] & (carry_g[DATA_WIDTH-2:1] & ~carry_d[DATA_WIDTH-3:0] 
 |  carry_d[DATA_WIDTH-2:1] & ~carry_g[DATA_WIDTH-3:0])
 | ~carry_p[DATA_WIDTH-1:2] & (carry_g[DATA_WIDTH-2:1] & ~carry_g[DATA_WIDTH-3:0] 
 |  carry_d[DATA_WIDTH-2:1] & ~carry_d[DATA_WIDTH-3:0]);


//==========================================================
//                     LZA coding
//==========================================================
assign data_for_ff1[DATA_WIDTH-1:0] = lza_precod[DATA_WIDTH-1:0] | upper_limit[DATA_WIDTH-1:0];
// &CombBeg; @66
always @( data_for_ff1[52:0])
begin
casez(data_for_ff1[DATA_WIDTH-1:0])
   53'b1????????????????????????????????????????????????????:lza_result[6:0] = 7'd0;
   53'b01???????????????????????????????????????????????????:lza_result[6:0] = 7'd1;
   53'b001??????????????????????????????????????????????????:lza_result[6:0] = 7'd2;
   53'b0001?????????????????????????????????????????????????:lza_result[6:0] = 7'd3;
   53'b00001????????????????????????????????????????????????:lza_result[6:0] = 7'd4;
   53'b000001???????????????????????????????????????????????:lza_result[6:0] = 7'd5;
   53'b0000001??????????????????????????????????????????????:lza_result[6:0] = 7'd6;
   53'b00000001?????????????????????????????????????????????:lza_result[6:0] = 7'd7;
   53'b000000001????????????????????????????????????????????:lza_result[6:0] = 7'd8;
   53'b0000000001???????????????????????????????????????????:lza_result[6:0] = 7'd9;
   53'b00000000001??????????????????????????????????????????:lza_result[6:0] = 7'd10;
   53'b000000000001?????????????????????????????????????????:lza_result[6:0] = 7'd11;
   53'b0000000000001????????????????????????????????????????:lza_result[6:0] = 7'd12;
   53'b00000000000001???????????????????????????????????????:lza_result[6:0] = 7'd13;
   53'b000000000000001??????????????????????????????????????:lza_result[6:0] = 7'd14;
   53'b0000000000000001?????????????????????????????????????:lza_result[6:0] = 7'd15;
   53'b00000000000000001????????????????????????????????????:lza_result[6:0] = 7'd16;
   53'b000000000000000001???????????????????????????????????:lza_result[6:0] = 7'd17;
   53'b0000000000000000001??????????????????????????????????:lza_result[6:0] = 7'd18;
   53'b00000000000000000001?????????????????????????????????:lza_result[6:0] = 7'd19;
   53'b000000000000000000001????????????????????????????????:lza_result[6:0] = 7'd20;
   53'b0000000000000000000001???????????????????????????????:lza_result[6:0] = 7'd21;
   53'b00000000000000000000001??????????????????????????????:lza_result[6:0] = 7'd22;
   53'b000000000000000000000001?????????????????????????????:lza_result[6:0] = 7'd23;
   53'b0000000000000000000000001????????????????????????????:lza_result[6:0] = 7'd24;
   53'b00000000000000000000000001???????????????????????????:lza_result[6:0] = 7'd25;
   53'b000000000000000000000000001??????????????????????????:lza_result[6:0] = 7'd26;
   53'b0000000000000000000000000001?????????????????????????:lza_result[6:0] = 7'd27;
   53'b00000000000000000000000000001????????????????????????:lza_result[6:0] = 7'd28;
   53'b000000000000000000000000000001???????????????????????:lza_result[6:0] = 7'd29;
   53'b0000000000000000000000000000001??????????????????????:lza_result[6:0] = 7'd30;
   53'b00000000000000000000000000000001?????????????????????:lza_result[6:0] = 7'd31;
   53'b000000000000000000000000000000001????????????????????:lza_result[6:0] = 7'd32;
   53'b0000000000000000000000000000000001???????????????????:lza_result[6:0] = 7'd33;
   53'b00000000000000000000000000000000001??????????????????:lza_result[6:0] = 7'd34;
   53'b000000000000000000000000000000000001?????????????????:lza_result[6:0] = 7'd35;
   53'b0000000000000000000000000000000000001????????????????:lza_result[6:0] = 7'd36;
   53'b00000000000000000000000000000000000001???????????????:lza_result[6:0] = 7'd37;
   53'b000000000000000000000000000000000000001??????????????:lza_result[6:0] = 7'd38;
   53'b0000000000000000000000000000000000000001?????????????:lza_result[6:0] = 7'd39;
   53'b00000000000000000000000000000000000000001????????????:lza_result[6:0] = 7'd40;
   53'b000000000000000000000000000000000000000001???????????:lza_result[6:0] = 7'd41;
   53'b0000000000000000000000000000000000000000001??????????:lza_result[6:0] = 7'd42;
   53'b00000000000000000000000000000000000000000001?????????:lza_result[6:0] = 7'd43;
   53'b000000000000000000000000000000000000000000001????????:lza_result[6:0] = 7'd44;
   53'b0000000000000000000000000000000000000000000001???????:lza_result[6:0] = 7'd45;
   53'b00000000000000000000000000000000000000000000001??????:lza_result[6:0] = 7'd46;
   53'b000000000000000000000000000000000000000000000001?????:lza_result[6:0] = 7'd47;
   53'b0000000000000000000000000000000000000000000000001????:lza_result[6:0] = 7'd48;
   53'b00000000000000000000000000000000000000000000000001???:lza_result[6:0] = 7'd49;
   53'b000000000000000000000000000000000000000000000000001??:lza_result[6:0] = 7'd50;
   53'b0000000000000000000000000000000000000000000000000001?:lza_result[6:0] = 7'd51;
   53'b00000000000000000000000000000000000000000000000000001:lza_result[6:0] = 7'd52;
   53'b00000000000000000000000000000000000000000000000000000:lza_result[6:0] = 7'd53;
  default                                                   :lza_result[6:0] = 7'd0;
endcase
// &CombEnd; @124
end

// &ModuleEnd; @126
endmodule


